module noDchu (
    input clk,D,ret,
    output reg q
);
  always @(posedge clk) begin
      
  end  
endmodule