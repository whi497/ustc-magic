module check (
    input clk,button,
    input [2:0] sw,
    output [4:0] out,[4:0] outin,[15:0] outstate
);
    parameter A = 4'ha;
    parameter B = 4'hb;
    parameter C = 4'hc;
    parameter D = 4'hd;
    wire [2:0] selsct;
endmodule